`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:09:01 12/01/2015 
// Design Name: 
// Module Name:    vgacontroller 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module vgacontroller(
    input resetbutton,
    input clk,
    output VGA_RED,
    output VGA_GREEN,
    output VGA_BLUE,
    output VGA_HSYNC,
    output VGA_VSYNC
    );

	//mod-2 counter
	reg mod2_reg;
	wire mod2_next;
	wire p_tick;
	//sync counters
	reg[9:0] h_count_reg, h_count_next;
	reg[9:0] v_count_reg, v_count_next;
	//output buffer
	reg v_sync_reg,h_sync_reg;
	wire v_sync_next,h_sync_next;
	//status signal
	wire h_end,v_end,pixel_tick;
	wire h_video_on,v_video_on,video_on;
	//pixels
	wire [9:0] pixel_x , pixel_y;
	//address
	reg [13:0] address=14'b00000000000000;
	//address counter
	wire [2:0] address_counter_next;
	reg [2:0] address_counter=3'b000;
//  RAMB16_S1  : In order to incorporate this function into the design,
//   Verilog   : the forllowing instance declaration needs to be placed
//  instance   : in the body of the design code.  The instance name
// declaration : (RAMB16_S1_inst) and/or the port declarations within the
//    code     : parenthesis may be changed to properly reference and
//             : connect this function to the design.  All inputs
//             : and outputs must be connected.

//  <-----Cut code below this line---->

   // RAMB16_S1: 16kx1 Single-Port RAM
   //            Spartan-3
   // Xilinx HDL Language Template, version 14.1

   RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
		//1bit to 4 , kathe init ine 2 grammes
      .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      // Address 4096 to 8191
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 12288 to 16383
      .INIT_30(256'h44444444444444444444444444444444FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_31(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_32(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_33(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_34(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_35(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_36(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_37(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_38(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_39(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3A(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3B(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3C(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3D(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3E(256'h4444444444444444444444444444444444444444444444444444444444444444),
      .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF44444444444444444444444444444444)
   ) RAMB16_S1_inst (
      .DO(VGA_RED),      // 1-bit Data Output
      .ADDR(address),  // 14-bit Address Input
      .CLK(p_tick),    // Clock
      .DI(1'b0),      // 1-bit Data Input
      .EN(1'b1),      // RAM Enable Input
      .SSR(1'b0),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );

  // End of RAMB16_S1_inst instantiation
//  RAMB16_S1  : In order to incorporate this function into the design,
//   Verilog   : the forllowing instance declaration needs to be placed
//  instance   : in the body of the design code.  The instance name
// declaration : (RAMB16_S1_inst) and/or the port declarations within the
//    code     : parenthesis may be changed to properly reference and
//             : connect this function to the design.  All inputs
//             : and outputs must be connected.

//  <-----Cut code below this line---->

   // RAMB16_S1: 16kx1 Single-Port RAM
   //            Spartan-3
   // Xilinx HDL Language Template, version 14.1

   RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
		//1bit to 4 , kathe init ine 2 grammes, kathe grammi 4x64=256 bits x16 ==> 4096
		//gia to aspro 4->c , 2->a , 1 ->9
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 4096 to 8191
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_21(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_22(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_23(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_24(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_25(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_26(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_27(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_28(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_29(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_2F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 12288 to 16383
      .INIT_30(256'h22222222222222222222222222222222FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_31(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_32(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_33(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_34(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_35(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_36(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_37(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_38(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_39(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3A(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3B(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3C(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3D(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3E(256'h2222222222222222222222222222222222222222222222222222222222222222),
      .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF22222222222222222222222222222222)	
   ) RAMB16_S3_inst (
      .DO(VGA_GREEN),      // 1-bit Data Output
      .ADDR(address),  // 14-bit Address Input
      .CLK(p_tick),    // Clock
      .DI(1'b0),      // 1-bit Data Input
      .EN(1'b1),      // RAM Enable Input
      .SSR(1'b0),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );

  // End of RAMB16_S1_inst instantiation
//  RAMB16_S1  : In order to incorporate this function into the design,
//   Verilog   : the forllowing instance declaration needs to be placed
//  instance   : in the body of the design code.  The instance name
// declaration : (RAMB16_S1_inst) and/or the port declarations within the
//    code     : parenthesis may be changed to properly reference and
//             : connect this function to the design.  All inputs
//             : and outputs must be connected.

//  <-----Cut code below this line---->

   // RAMB16_S1: 16kx1 Single-Port RAM
   //            Spartan-3
   // Xilinx HDL Language Template, version 14.1

   RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("WRITE_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
		//1bit to 4 , kathe init ine 2 grammes
      .INIT_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_0F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 4096 to 8191
      .INIT_10(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_11(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_12(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_13(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_14(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_15(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_16(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_17(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_18(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_19(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1A(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1B(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1C(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1D(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1E(256'h0000000000000000000000000000000000000000000000000000000000000000),
      .INIT_1F(256'h0000000000000000000000000000000000000000000000000000000000000000),
      // Address 8192 to 12287
      .INIT_20(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_24(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_25(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_26(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_27(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_28(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_29(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_2A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_2B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_2C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_2D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_2E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      .INIT_2F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000000000000000000000000),
      // Address 12288 to 16383
      .INIT_30(256'h11111111111111111111111111111111FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_31(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_32(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_33(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_34(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_35(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_36(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_37(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_38(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_39(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3A(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3B(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3C(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3D(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3E(256'h1111111111111111111111111111111111111111111111111111111111111111),
      .INIT_3F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF11111111111111111111111111111111)
   ) RAMB16_BLUE_inst (
      .DO(VGA_BLUE),      // 1-bit Data Output
      .ADDR(address),  // 14-bit Address Input
      .CLK(p_tick),    // Clock
      .DI(1'b0),      // 1-bit Data Input
      .EN(1'b1),      // RAM Enable Input
      .SSR(1'b0),    // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );

  // End of RAMB16_S1_inst instantiation  
//contant declartion
// VGA 640x480 parameters	
	localparam HD =640; // horizontal display area
	localparam HF =48;  // h.front (left) border
	localparam HB =16;  // h. back (right) border
	localparam HR =96;  // h.retrace
	localparam VD =480; // vertical display area
	localparam VF =10;  // v.front(top) border
	localparam VB =33;  // v.back (bottom) border
	localparam VR =2;   // v.retace


	always @(posedge clk,posedge resetbutton)
		if(resetbutton)
			begin
				mod2_reg <= 1'b0;
				v_count_reg <= 0;
				h_count_reg <= 0;
				v_sync_reg <= 1'b0;
				h_sync_reg <= 1'b0;
				//address_counter <= 1'b0;	
			end
		else
			begin
				mod2_reg <= mod2_next;
				v_count_reg <= v_count_next;
				h_count_reg <= h_count_next;
				v_sync_reg <= v_sync_next;
				h_sync_reg <= h_sync_next;
				//address_counter <= address_counter_next;
			end
	
	
	//mod-2 circuit to generate 25 Mhz enable tick
	assign mod2_next = ~mod2_reg;
	assign pixel_tick = mod2_reg;
	//end of horizontial counter (799)
	assign h_end = ( h_count_reg == ( HD + HF + HB + HR -2));
	
	//end of vertical counter (524)
	assign v_end =( v_count_reg == ( VD + VF + VB + VR -1));

	//assign address_counter_next = address_counter + 1;
	// next-state logic of mod-800 horizontal sync coumter
	always @(clk)
		if(pixel_tick)
			if( h_end)
				h_count_next = 0;
			else
				h_count_next = h_count_reg + 1;
		else
			h_count_next = h_count_reg;
			
	// next-state logic of mod-525 vertical sunc counter
	always @(clk)
		if(pixel_tick & h_end)
			if(v_end)
				v_count_next <= 0;
			else 
				v_count_next <= v_count_reg + 1;
		else
			v_count_next <= v_count_reg;
	

	always@(pixel_tick)
		if( address_counter == 5) //dn me afine mod 5
			begin
			address <= address +1;
			address_counter <= 0;
			end
		else 
			address_counter <= address_counter + 1;
	
	
	
	//horizontal and vertical sync buffered
	//h_sync_nect asserted between 656 and 751
	
	assign h_sync_next = (h_count_reg >= (HD+HB-1) && h_count_reg <= (HD+HB+HR-2));
	
	//v_sync_nect asserted between 490 and 491
	
	assign v_sync_next = (v_count_reg >= ((VD+VF-1)) && v_count_reg <= (VD+VF ));
	
	//address ++ when pixel_x % 5 == 0
	
	//assign address = ((pixel_x % 5) == 0 ) ? (address+1): (address); 

	//video enable
	assign h_video_on = ((h_count_reg < HD )) ; 
	assign v_video_on = (v_count_reg < VD ) ;

	//output
	assign VGA_HSYNC = h_sync_reg;
	assign VGA_VSYNC = v_sync_reg;
	assign pixel_x = h_count_reg;
	assign pixel_y = v_count_reg;
	assign p_tick = pixel_tick;

endmodule
